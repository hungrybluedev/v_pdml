module spec

pub struct PMLTestSuite {
pub:
	name  string
	desc  string
	cases []PMLTestCase
}
