module pml
